module shift(


);

endmodule
