module incrementR (
	input inc,
	input reset_n,
	input clk50,
	output [7:0] value,
	output reg [romsize-1:0] Iaddress

	
);

parameter romsize = 14;

//output reg [romsize-1:0] Iaddress;





endmodule
